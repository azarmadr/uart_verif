typedef enum{
	MEM	=0,
	REG	=1} mem_reg_t;
typedef enum{
	READ	=0,
	WRITE	=1} wr_rd_t;

